VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ws_ip__logo
  CLASS BLOCK ;
  FOREIGN gf180mcu_ws_ip__logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 400 BY 400 ;
  OBS
      LAYER Metal5 ;
        RECT 0.0 0.0 400 400 ;
  END
END gf180mcu_ws_ip__logo
END LIBRARY

