module gf180mcu_ws_ip__ce_logo;
endmodule
